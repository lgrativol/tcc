library ieee;
use ieee.std_logic_1164.all;

package sim_input_pkg is
   constant SIM_INPUT_TARGETFREQ     : positive  := 100000;
   constant SIM_INPUT_NBCYCLES       : natural   := 200;
end sim_input_pkg;
